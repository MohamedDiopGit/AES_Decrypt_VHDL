library IEEE;
use IEEE.std_logic_1164.all;

library LIB_AES;
use LIB_AES.state_definition_package.all;

configuration InvShiftRows_conf of InvShiftRows is
	for InvShiftRows_arch-- architecture name
	end for;
end InvShiftRows_conf;
