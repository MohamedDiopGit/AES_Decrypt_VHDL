library IEEE;
use IEEE.std_logic_1164.all;

library LIB_RTL;


configuration AddRoundKey_conf of AddRoundKey is
	for AddRoundKey_arch-- architecture name
	end for;
end AddRoundKey_conf;
