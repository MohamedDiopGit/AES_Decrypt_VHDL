library IEEE;
use IEEE.std_logic_1164.all;

library LIB_AES;
use LIB_AES.state_definition_package.all;

configuration InvMixColumnsX_conf of InvMixColumnsX is
	for InvMixColumnsX_arch -- architecture name
	end for;
end InvMixColumnsX_conf;
